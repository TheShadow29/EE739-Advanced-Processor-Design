library ieee ;
use ieee.std_logic_1164.all ;
library work;

package dispatch_components is
	
end package;