library ieee ;
use ieee.std_logic_1164.all ;
library work;

package writeback_components is
end package;